`ifndef _
`define _

//TODO Module 
//
// 
//
module ;
endmodule

`endif
