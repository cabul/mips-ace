`ifndef _icache
`define _icache

//////////////////////
// Instruction Cache
//
module icache;
endmodule

`endif
