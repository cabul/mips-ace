`include "alu.v"

module alu_tb;

initial begin
	$monitor("Success.");
end

endmodule;