`ifndef _dcache
`define _dcache

//TODO Module dcache
///
/// dcache
///
module dcache;
endmodule

`endif
